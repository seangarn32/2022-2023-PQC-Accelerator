library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.globals.all;

entity processing_element_i is
    port (
        
        A   : in    standard_
    );
end entity;

architecture rtl of processing_element_i is
end architecture;