library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.globals.all;

entity pqc_accelerator_top is
end entity;

architecture rtl of pqc_accelerator_top is
end architecture;