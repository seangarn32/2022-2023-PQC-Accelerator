library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.globals_pkg.all;

entity fsm is
    port ( 
        reset : in  STD_LOGIC;
        start : in  STD_LOGIC;
        clk : in  STD_LOGIC
    );
end fsm;

architecture rtl of fsm is

    type state_available is (SETUP, DATA_IN, PE, DATA_OUT);  --type of state machine.
    signal present_state,next_state: state_available;
    signal counter: STD_LOGIC_VECTOR(7 downto 0);
    signal counter_ena: STD_LOGIC;
    signal counter_reset: STD_LOGIC;

begin
    process (clk,reset)
    begin
        if (reset='1') then
            present_state<= SETUP;  --default state on reset.
        elsif (rising_edge(clk)) then
            present_state<= next_state;   --state change.
        end if;
    end process;

    STATE_COUNTER: entity work.counter(rtl)
            port map (
                clk, counter_reset, counter_ena, counter
            );

    process (present_state)
    begin
        case present_state is
            when SETUP =>        --when current state is "A"
                counter_reset <= '1';
                if(start ='0') then
                    next_state <= SETUP;
                else
                    next_state <= DATA_IN; -- once we flip a switch, it will move to DATA_IN
                end if;  
            when DATA_IN =>        --when current state is "B"
                counter_ena <= '1';
                if(counter > "00010000") then
                    next_state <= PE;
                    counter_ena <= '0';
                else
                    next_state<= DATA_IN;
                end if;
            when PE =>       --when current state is "C"
                counter_ena <= '1';
                if(counter = "11111111") then
                    next_state <= DATA_OUT;
                    counter_ena <= '0';
                else
                    next_state<= PE;
                end if;
            when DATA_OUT =>         --when current state is "D"
                counter_ena <= '1';
                if(counter = "11111111") then
                    next_state <= SETUP;
                    counter_ena <= '0';
                else
                    next_state<= DATA_OUT;
                end if;
        end case;
    end process;
end rtl;
