library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package globals_pkg is

    constant N_SIZE : integer := 8;

end package;